module alu_control(control_signal);